
    module KEY_OR_LED ( A, B, F );
        input A, B;         // ??????
        output F;           // ??????
        assign F = A||B;    //??F??1 LED?????
                            //??F??0 LED????
    endmodule
