
module SMG_LED (led_bit,dataout);

//input clk_50M ;       //????50M?? ?17????
output [7:0] dataout;   //????????ABCDEFG????????????
output led_bit;         //?????????

reg [7:0] dataout;
reg       led_bit;  

//always @ ( posedge clk_50M )

 //begin
 always  led_bit <= 'b0; //??????????????

 always  dataout<=8'b11000000; //??7????????????
                               //?????????0?9?????A?F,????????????
                               //????????????0

 //end
endmodule

