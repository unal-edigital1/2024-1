
    module KEY_NAND_LED ( A,B,F );
    input A,B;            // ??????
    output F;             // ??????
    assign F =~(A & B);   //??A B???1 ;LED?????
                          //??A B??????? LED????
    endmodule
