

module ledwater (clk_50M,led_out);
input   clk_50M;       //??????50M  input  pin17
                       //????????50,000,000HZ

output  led_out;       //???????

reg [24:0] count;  //??????25,000,000HZ
reg  div_clk;     //??????????????????
reg  led_out;

//?????????????
always @ ( posedge clk_50M )
begin
if ( count==25000000 )
 begin     //??????????????50,000,000HZ
           //?????count??????????25,000,000HZ
  div_clk<=~div_clk;  //?????????0.5?????????
                      //????????1Hz??????
   count<=0;          //???????
  end
else
  count<=count+1;     //??????
  led_out <= div_clk;  //??????????????????
                      //?LED????????
end 

endmodule














